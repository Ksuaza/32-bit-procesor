library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

entity Salidas is port (
 Data :in std_logic_vector (31 downto 0);
 Direccion :in std_logic_vector (2 downto 0);
 W :in std_logic
);
end Salidas;

architecture interna of Salidas is
begin

end interna;

--Kevin Suaza