library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

entity Entradas is port (
Q :out std_logic_vector (31 downto 0)
);
end Entradas;

architecture interna of Entradas is
begin

end interna;

--Kevin Suaza